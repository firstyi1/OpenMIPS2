`include "defines.v"

module mem(
    input   wire                rst     ,

    // 来自exe阶段的信息
    input   wire [`RegAddrBus]  wd_i    ,
    input   wire                wreg_i  ,
    input   wire [`RegBus]      wdata_i ,

    // mem阶段的结果
    output  reg  [`RegAddrBus]  wd_o    ,
    output  reg                 wreg_o  ,
    output  reg [`RegBus]       wdata_o

);

    // 目前只实现了 ori 指令，且该指令没有mem阶段，因此当前mem阶段不进行操作
    always @(*) begin
        if (rst == `RstEnable) begin
            wd_o    <= `NOPRegAddr;
            wreg_o  <= `WriteDisable;
            wdata_o <= `ZeroWord;
        end
        else begin
            wd_o    <= wd_i;
            wreg_o  <= wreg_i;
            wdata_o <= wdata_i;
        end
    end

endmodule